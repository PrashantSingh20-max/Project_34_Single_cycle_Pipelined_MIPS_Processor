
//comparator comp(equala,equalb,equalD);
module comparator(
		  input [5:0]a,b,
		  output c

);

assign c=(a==b);
endmodule